--------------------------------------------------------------------------------
-- PICT MEM
-- Anders Nilsson
-- 16-feb-2016
-- Version 1.1


-- library declaration
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;            -- basic IEEE library
use IEEE.NUMERIC_STD.ALL;               -- IEEE library for the unsigned type


-- entity
entity PICT_MEM is
  port ( clk		: in std_logic;
         -- port 1;
         --addr1		: in unsigned(10 downto 0);
         -- port 2
         data_out2	: out std_logic_vector(3 downto 0);
         addr2		: in unsigned(12 downto 0));

end PICT_MEM;

	
-- architecture
architecture Behavioral of PICT_MEM is

  -- picture memory type
  type ram_t is array (0 to 4799) of std_logic_vector(3 downto 0);
  -- initiate picture memory to one cursor ("1F") followed by spaces ("00")
  signal pictMem : ram_t := (
x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"2",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"2",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"2",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"2",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"2",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"2",x"2",x"2",x"2",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"1",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"5",x"0", 
 
x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
);


begin

  process(clk)
  begin
    if rising_edge(clk) then
      data_out2 <= pictMem(to_integer(addr2));
    end if;
  end process;


end Behavioral;

