library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- uMem interface
entity uMem is
  port (
    uAddr : in unsigned(7 downto 0);
    uData : out unsigned(24 downto 0));
end uMem;

architecture Behavioral of uMem is

-- micro Memory
type u_mem_t is array (0 to 90) of unsigned(24 downto 0);
constant u_mem_c : u_mem_t :=
   --ALU__TB__FB_PC_LC_SEQ__uAddr
  (b"0000_011_111_0_00_0000_00000000",   --ASR := PC
   b"0000_010_001_1_00_0000_00000000",   --IR := PM , PC := PC+1
   b"0000_000_000_0_00_0010_00000000",   -- uPC := K2(Mod) 
   b"0000_010_110_0_00_0000_00000000",   -- Grx := PM(A) LOAD 
   b"0000_000_000_0_00_0011_00000000",   
   b"0000_000_000_0_00_1111_00000000",   --HALT undone
   b"0000_000_000_0_00_0011_00000000",
   b"0000_110_010_0_00_0000_00000000",   --STORE
   b"0000_000_000_0_00_0011_00000000",
   b"0001_110_000_0_00_0000_00000000",   --ADD
   b"0100_010_000_0_00_0000_00000000",
   b"0000_100_110_0_00_0000_00000000",
   b"0000_000_000_0_00_0011_00000000",
   b"0001_110_000_0_00_0000_00000000",   --SUB
   b"0101_010_000_0_00_0000_00000000",
   b"0000_100_110_0_00_0000_00000000",
   b"0000_000_000_0_00_0011_00000000",
   b"0001_110_000_0_00_0000_00000000",   --AND
   b"0110_010_000_0_00_0000_00000000",
   b"0000_100_110_0_00_0000_00000000",
   b"0000_000_000_0_00_0011_00000000",
   b"0000_010_011_0_00_0000_00000000",  -- BRA
   b"0000_000_000_0_00_0011_00000000",
   b"0001_110_000_0_00_0000_00000000",  -- CMP
   b"0101_010_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0011_00000000",
   b"0000_000_000_0_00_1000_00010101",  -- BEQ
   b"0000_000_000_0_00_0011_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0011_00000000",
   b"0000_000_000_0_00_1001_00100001",  --BGE
   b"0000_000_000_0_00_1011_00100010",
   b"0000_000_000_0_00_0101_00010101",
   b"0000_000_000_0_00_1011_00100011",
   b"0000_000_000_0_00_0011_00000000",
   b"0000_000_000_0_00_0101_00010101",
   b"0001_110_000_0_00_0000_00000000",  -- MULU
   b"0000_010_000_0_10_0000_00000000", 
   b"0000_000_000_0_00_1100_00101001",
   b"0100_110_000_0_01_0000_00000000",
   b"0000_000_000_0_00_0101_00100110",
   b"0000_100_110_0_00_0000_00000000",
   b"0000_000_000_0_00_0011_00000000",
   b"0000_001_111_0_00_0001_00000000",  -- Direct
   b"0000_001_111_0_00_0000_00000000",  -- Indirect
   b"0000_010_111_0_00_0001_00000000",
   b"0000_011_111_1_00_0001_00000000",  -- immediate
   b"0000_000_000_0_00_0011_00000000",  
   b"0000_010_111_0_00_0000_00000000",  --Tra
   b"1100_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0011_00000000",
   b"0001_011_000_0_00_0000_00000000",  -- BRA_PLUS
   b"0100_010_000_0_00_0000_00000000",
   b"0000_100_011_0_00_0000_00000000",
   b"0000_000_000_0_00_0011_00000000",
   b"0001_011_000_0_00_0000_00000000",  -- BRA_MINUS
   b"0101_010_000_0_00_0000_00000000",
   b"0000_100_011_0_00_0000_00000000",
   b"0000_000_000_0_00_0011_00000000",
   b"0000_000_000_0_00_0101_00111000",
   b"0000_000_000_0_00_0011_00000000",
   b"0000_000_000_0_00_1000_00111111",  -- BNE
   b"0000_000_000_0_00_0101_00010101",
   b"0000_000_000_0_00_0011_00000000",
   b"0000_000_000_0_00_1001_01000011",  --BL 40
   b"0000_000_000_0_00_1011_01000100",
   b"0000_000_000_0_00_0011_00000000",
   b"0000_000_000_0_00_1011_01000010",
   b"0000_000_000_0_00_0101_00010101",
   b"1110_000_000_0_11_0000_11111111",  --BEEP
   b"0000_000_000_0_00_1100_01001000",
   b"0000_000_000_0_01_0000_01000110",
   b"1111_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0011_00000000",
   b"0000_001_111_0_00_0000_00000000",  --Inception
   b"0000_010_111_0_00_0000_00000000",
   b"0000_010_111_0_00_0001_00000000",
   b"0000_000_000_0_00_0011_00000000",
   others =>(others => '0'));

signal u_mem : u_mem_t := u_mem_c;

begin  -- Behavioral
  uData <= u_mem(to_integer(uAddr));

end Behavioral;
