library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- uMem interface
entity uMem is
  port (
    uAddr : in unsigned(7 downto 0);
    uData : out unsigned(24 downto 0));
end uMem;

architecture Behavioral of uMem is

-- micro Memory
type u_mem_t is array (0 to 39) of unsigned(24 downto 0);
constant u_mem_c : u_mem_t :=
   --ALU__TB__FB_PC_LC_SEQ__uAddr
  (b"0000_011_111_0_00_0000_00000000",   --ASR := PC
   b"0000_010_001_1_00_0000_00000000",   --IR := PM , PC := PC+1
   b"0000_001_111_0_00_0001_00000000",   -- ASR := IR , uPC := K1 
   b"0000_010_110_0_00_0000_00000000",   -- Grx := PM(A) LOAD
   b"0000_000_000_0_00_0011_00000000",   
   b"0000_000_000_0_00_1111_00000000",   --HALT
   b"0000_000_000_0_00_0011_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000",
   b"0000_000_000_0_00_0000_00000000");

signal u_mem : u_mem_t := u_mem_c;

begin  -- Behavioral
  uData <= u_mem(to_integer(uAddr));

end Behavioral;
