library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

--CPU interface
entity proj is
  port(clk: in std_logic;
       rst: in std_logic;
       tile: out unsigned(3 downto 0);
       index: out unsigned(15 downto 0));
end proj ;

architecture Behavioral of proj is


  -- micro Memory component
  component uMem
    port(uAddr : in unsigned(7 downto 0);
         uData : out unsigned(24 downto 0));
  end component;

  -- program Memory component
 -- component pMem
   -- port(pAddr : in unsigned(31 downto 0);
     --    pData : out unsigned(31 downto 0));
 -- end component;
  

  
  -- K1 memory component
  component K1
    port(operand: in unsigned(3 downto 0);
         K1_adress: out unsigned(7 downto 0));
  end component;

   -- K1 memory component
  component K2
    port(modd: in unsigned(3 downto 0);
         K2_adress: out unsigned(7 downto 0));
  end component;

  --K2 memory component
  signal K2_reg : unsigned(7 downto 0); --K2 memory output
  -- K1 memory component
  signal K1_reg : unsigned(7 downto 0);  -- K1 memory output
  -- micro memory signals
  signal uM : unsigned(24 downto 0); -- micro Memory output
  signal uPC : unsigned(7 downto 0); -- micro Program Counter
  --signal uPCsig : std_logic; -- (0:uPC++, 1:uPC=uAddr)
  signal uAddr : unsigned(7 downto 0); -- micro Address
  signal TB : unsigned(2 downto 0); -- To Bus field
  signal FB : unsigned(2 downto 0); -- From Bus field
  signal ALU : unsigned(3 downto 0); -- ALU for arithmetical/logical operations
  signal LC : unsigned(1 downto 0) ; -- loop counter
  signal SEQ : unsigned(3 downto 0); -- uPC contidion setter

  -- program memory signals
  signal PM : unsigned(31 downto 0); -- Program Memory output
  signal PC : unsigned(31 downto 0); -- Program Counter
  signal Pcsig : std_logic; -- 0:PC=PC, 1:PC++
  signal ASR : unsigned(31 downto 0); -- Address Register
  signal IR : unsigned(31 downto 0); -- Instruction Register
  signal DATA_BUS : unsigned(31 downto 0); -- Data Bus
  signal AR : unsigned(32 downto 0) := ('0' & x"00000000"); -- stores alu operated values
  signal GRx : unsigned(3 downto 0) ; -- grx part in pm
  signal OP : unsigned(3 downto 0); -- Oeration part in pm
  signal GRx0 : unsigned(31 downto 0); 		
  signal GRx1 : unsigned(31 downto 0); 	
  signal GRx2 : unsigned(31 downto 0); 	
  signal GRx3 : unsigned(31 downto 0); 	
  signal LC_REG : unsigned(15 downto 0):= x"0000"; -- register holding loop value
  signal L , N, Z, O, C : std_logic := '0';    -- flags
  signal HALT : std_logic := '1';       -- flag for halting PC
  signal PM_ADR : unsigned(15 downto 0);  -- adress part of PM
  signal AR_TEMP : std_logic :='0';  -- temporary value for MSB in AR
  signal ADR_MOD : unsigned(3 downto 0);  -- Adress mod part of PM
  --signal index : unsigned(15 downto 0) := x"0000";  -- index for pict_mem
  signal indexbuffer : unsigned(15 downto 0) := "1111111111111111";  -- index buffer

  -----------------------------------------------------------------------------
  -- PRIMARY MEMMORY
  -----------------------------------------------------------------------------
  type p_mem_t is array (0 to 5000) of unsigned(31 downto 0);
  constant p_mem_c : p_mem_t :=
    (x"00200000",                       -- load 2 till GR0
     x"00000002",                       
     x"20000019",                       -- store Gr0 i $1B
     x"00200000",                       -- load 3000 till gr0
     x"00000BB8",
     x"40200000",                      
     x"00000001",                       -- 1 till gr0
     x"B000000C",
     x"70200000",                       -- CMP gr0 och 1
     x"00000001",
     x"9000000B",                       -- BGE hoppa till $05
     x"00000005",
     x"00000019",
     x"10000000",
     x"00000000",
     x"00000000",
     x"00000000",
     x"00000000",
     x"00000000",
     x"00000000",
     x"00000000",
     x"00000000",
     x"00000000",
     x"00000000",
     x"00000000",
     x"00000000",
     x"60000006",                       --1A


     others => (others => '0'));

  signal p_mem : p_mem_t := p_mem_c;


-------------------------------------------------------------------------------
-- --------------------------------------------------------------------------
-------------------------------------------------------------------------------











  
begin

  
  -- mPC : micro Program Counter
  process(clk)
  begin
    if rising_edge(clk) then
      if (rst = '1' or SEQ = "0011") then
        uPC <= (others => '0');
      elsif (SEQ ="0101") then
        uPC <= uAddr;
      elsif (SEQ = "0000") then
        uPC <= uPC + 1;
      elsif (SEQ="0001") then
        uPC <= K1_reg;
      elsif (SEQ = "0010") then
        uPC <= K2_reg;
      elsif (SEQ = "1000" and Z='1') then
        uPC <= uAddr;
      elsif (SEQ = "1001" and N='1') then
        uPC <= uAddr;
      elsif (SEQ = "1100" and L='1') then
        uPC <= uAddr;
      elsif (SEQ ="1010" and C = '1') then
        uPC <= uAddr;
      elsif (SEQ="1011" and O = '1') then
        uPC <= uAddr;
      elsif (SEQ = "1111") then
        HALT <= '0';
      else
        uPC <= uPC + 1;
      end if;
    end if;
  end process;
	
  -- PC : Program Counter
  process(clk)
  begin
    if (HALT ='1') then  
      if rising_edge(clk) then
        if (rst = '1') then
          PC <= (others => '0');
        elsif (FB = "011") then
          PC <= DATA_BUS;
        elsif (PCsig = '1') then
          PC <= PC + 1;
        end if;
      end if;
    end if;
  end process;
	
  -- IR : Instruction Register
  process(clk)
  begin
    if rising_edge(clk) then
      if (rst = '1') then
        IR <= (others => '0');
      elsif (FB = "001") then
        IR <= DATA_BUS;
      end if;
    end if;
  end pRocess;
	
  -- ASR : Address Register
  process(clk)
  begin
    if rising_edge(clk) then
      if (rst = '1') then
        ASR <= (others => '0');
      elsif (FB = "111") then
        ASR <= x"0000" & DATA_BUS(15 downto 0);
       
     end if;
	
    end if;
  end process;

  -- PM
  process(clk)
  begin
    if rising_edge(clk) then
      if (FB ="010") then
        p_mem(to_integer(ASR)) <= DATA_BUS;
      
      end if;
    end if;
  end process;
  
  -- GRx: general register
  process(clk)
  begin
    if rising_edge(clk) then 
      if (rst ='1') then
	GRx0 <= (others => '0');
	GRx1 <= (others => '0');
	GRx2 <= (others => '0');
	GRx3 <= (others => '0');
      elsif (FB = "110") then
	if (GRx = 0) then
	   GRx0 <= DATA_BUS;
	elsif (GRx = 1) then
	   GRx1 <= DATA_BUS;
	elsif (GRx = 2) then
	   GRx2 <= DATA_BUS;
        elsif (GRx = 3) then
    	   GRx3 <= DATA_BUS;
	end if;
      end if;
    end if;
  end process;	
 


 --LC
 process(clk)
   begin
     if rising_edge(clk) then
       if (rst='1') then
         LC_REG <= (others => '0');
       elsif (LC = "01") then
         LC_REG <= LC_REG - 1;
       elsif (LC = "10") then
         LC_REG <= DATA_BUS(15 downto 0);
       elsif (LC ="11") then
         LC_REG <= x"00" & uAddr;
       end if;
     end if;
 end process;

 -- ALU  
 process(clk)
   
 begin
    if rising_edge(clk) then
      AR_TEMP <= AR(31);
      if (rst ='1' or ALU = "0011") then
        AR <= (others => '0');
      elsif (ALU= "0001") then
        AR <= ('0' & DATA_BUS);
        
      elsif (ALU ="0100") then
        AR <= AR + ('0' & DATA_BUS);
     
     
        
      Elsif (ALU ="0101") then
        AR <= AR - ('0' & DATA_BUS);
       
      elsif (ALU = "0110") then
        AR <= AR and ('0' & DATA_BUS);
          
      elsif (ALU = "0111") then
        AR <= AR or ('0' & DATA_BUS);

      elsif ( ALU = "1100") then
        tile <= PM(3 downto 0);
        indexbuffer <= indexbuffer +1;
        if (indexbuffer = 1) then
          indexbuffer <= (others => '0');
        end if;
        
      end if; 
    end if;
 end process;                           

  -- micro memory component connection
  U0 : uMem port map(uAddr=>uPC, uData=>uM);

  -- K2 memory component connection
  U1 : K2 port map (modd => ADR_MOD, K2_adress => K2_reg);
 

  -- K1 memory component connection
  U2 : K1 port map(operand => OP, K1_adress => K1_reg);


  -- Pict_mem index
  index <= indexbuffer;
     
  -- ALU Flags
    -- AR_TEMP <= AR(31);
     Z <= '1' when (AR = 0) else '0';
     N <= '1' when (signed(AR)<0) else '0';
     C <= '1' when (AR(32) = '1')  else '0';
     O <= '1' when ((AR(31)/=AR_TEMP) and (AR(31)= DATA_BUS(31))) else '0';
     L <= '1' when (LC_REG = 0) else '0';
  
  -- micro memory signal assignments
  
  uAddr <= uM(7 downto 0);
  SEQ <= uM(11 downto 8);
  LC <= uM(13 downto 12);
  PCsig <= uM(14);
  FB <= uM(17 downto 15);
  TB <= uM(20 downto 18);
  ALU <= uM(24 downto 21);       
  	
  -- primary memory signal assignment
 
  PM <= p_mem(to_integer(ASR));
  GRx <= IR(27 downto 24);
  OP <= IR(31 downto 28);
  PM_ADR <= IR(15 downto 0);
  ADR_MOD <= IR(23 downto 20);   
  -- data bus assignment
  DATA_BUS <= IR when (TB = "001") else
    PM when (TB = "010") else
    PC when (TB = "011") else
    AR(31 downto 0) when (TB = "100") else
    GRx0 when (TB ="110" and GRx = 0) else
    GRx1 when (TB ="110" and GRx = 1) else
    GRx2 when (TB ="110" and GRx = 2) else
    GRx3 when (TB ="110" and GRx = 3) else
    (others => '0');

end Behavioral;
